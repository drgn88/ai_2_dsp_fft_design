`timescale 1ns / 1ps

module twf_rom_mod12 #(
    parameter ROM_DEPTH = 512,
    parameter TWF_WIDTH = 9,
    parameter ADDR_WIDTH = 9,
    parameter OFFSET = 8
) (
    // input clk,
    input [ADDR_WIDTH-1:0] addr,
    //input en,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_R_add,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_Q_add,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_R_sub,
    output logic signed [TWF_WIDTH-1:0] twiddle_fac_Q_sub
);

    logic signed [TWF_WIDTH-1:0] rom_real_data[ROM_DEPTH-1:0];
    logic signed [TWF_WIDTH-1:0] rom_imag_data[ROM_DEPTH-1:0];

	assign twiddle_fac_R_add = rom_real_data[addr];
    assign twiddle_fac_Q_add = rom_imag_data[addr];
    assign twiddle_fac_R_sub = rom_real_data[addr+OFFSET];
    assign twiddle_fac_Q_sub = rom_imag_data[addr+OFFSET];


    assign rom_real_data[0]   = 128;
	assign rom_real_data[1]   = 128;
	assign rom_real_data[2]   = 128;
	assign rom_real_data[3]   = 128;
	assign rom_real_data[4]   = 128;
	assign rom_real_data[5]   = 128;
	assign rom_real_data[6]   = 128;
	assign rom_real_data[7]   = 128;
	assign rom_real_data[8]   = 128;
	assign rom_real_data[9]   = 118;
	assign rom_real_data[10]  = 91;
	assign rom_real_data[11]  = 49;
	assign rom_real_data[12]  = 0;
	assign rom_real_data[13]  = -49;
	assign rom_real_data[14]  = -91;
	assign rom_real_data[15]  = -118;
	assign rom_real_data[16]  = 128;
	assign rom_real_data[17]  = 126;
	assign rom_real_data[18]  = 118;
	assign rom_real_data[19]  = 106;
	assign rom_real_data[20]  = 91;
	assign rom_real_data[21]  = 71;
	assign rom_real_data[22]  = 49;
	assign rom_real_data[23]  = 25;
	assign rom_real_data[24]  = 128;
	assign rom_real_data[25]  = 106;
	assign rom_real_data[26]  = 49;
	assign rom_real_data[27]  = -25;
	assign rom_real_data[28]  = -91;
	assign rom_real_data[29]  = -126;
	assign rom_real_data[30]  = -118;
	assign rom_real_data[31]  = -71;
	assign rom_real_data[32]  = 128;
	assign rom_real_data[33]  = 127;
	assign rom_real_data[34]  = 126;
	assign rom_real_data[35]  = 122;
	assign rom_real_data[36]  = 118;
	assign rom_real_data[37]  = 113;
	assign rom_real_data[38]  = 106;
	assign rom_real_data[39]  = 99;
	assign rom_real_data[40]  = 128;
	assign rom_real_data[41]  = 113;
	assign rom_real_data[42]  = 71;
	assign rom_real_data[43]  = 13;
	assign rom_real_data[44]  = -49;
	assign rom_real_data[45]  = -99;
	assign rom_real_data[46]  = -126;
	assign rom_real_data[47]  = -122;
	assign rom_real_data[48]  = 128;
	assign rom_real_data[49]  = 122;
	assign rom_real_data[50]  = 106;
	assign rom_real_data[51]  = 81;
	assign rom_real_data[52]  = 49;
	assign rom_real_data[53]  = 13;
	assign rom_real_data[54]  = -25;
	assign rom_real_data[55]  = -60;
	assign rom_real_data[56]  = 128;
	assign rom_real_data[57]  = 99;
	assign rom_real_data[58]  = 25;
	assign rom_real_data[59]  = -60;
	assign rom_real_data[60]  = -118;
	assign rom_real_data[61]  = -122;
	assign rom_real_data[62]  = -71;
	assign rom_real_data[63]  = 13;
	assign rom_real_data[64]  = 128;
	assign rom_real_data[65]  = 128;
	assign rom_real_data[66]  = 128;
	assign rom_real_data[67]  = 128;
	assign rom_real_data[68]  = 128;
	assign rom_real_data[69]  = 128;
	assign rom_real_data[70]  = 128;
	assign rom_real_data[71]  = 128;
	assign rom_real_data[72]  = 128;
	assign rom_real_data[73]  = 118;
	assign rom_real_data[74]  = 91;
	assign rom_real_data[75]  = 49;
	assign rom_real_data[76]  = 0;
	assign rom_real_data[77]  = -49;
	assign rom_real_data[78]  = -91;
	assign rom_real_data[79]  = -118;
	assign rom_real_data[80]  = 128;
	assign rom_real_data[81]  = 126;
	assign rom_real_data[82]  = 118;
	assign rom_real_data[83]  = 106;
	assign rom_real_data[84]  = 91;
	assign rom_real_data[85]  = 71;
	assign rom_real_data[86]  = 49;
	assign rom_real_data[87]  = 25;
	assign rom_real_data[88]  = 128;
	assign rom_real_data[89]  = 106;
	assign rom_real_data[90]  = 49;
	assign rom_real_data[91]  = -25;
	assign rom_real_data[92]  = -91;
	assign rom_real_data[93]  = -126;
	assign rom_real_data[94]  = -118;
	assign rom_real_data[95]  = -71;
	assign rom_real_data[96]  = 128;
	assign rom_real_data[97]  = 127;
	assign rom_real_data[98]  = 126;
	assign rom_real_data[99]  = 122;
	assign rom_real_data[100] = 118;
	assign rom_real_data[101] = 113;
	assign rom_real_data[102] = 106;
	assign rom_real_data[103] = 99;
	assign rom_real_data[104] = 128;
	assign rom_real_data[105] = 113;
	assign rom_real_data[106] = 71;
	assign rom_real_data[107] = 13;
	assign rom_real_data[108] = -49;
	assign rom_real_data[109] = -99;
	assign rom_real_data[110] = -126;
	assign rom_real_data[111] = -122;
	assign rom_real_data[112] = 128;
	assign rom_real_data[113] = 122;
	assign rom_real_data[114] = 106;
	assign rom_real_data[115] = 81;
	assign rom_real_data[116] = 49;
	assign rom_real_data[117] = 13;
	assign rom_real_data[118] = -25;
	assign rom_real_data[119] = -60;
	assign rom_real_data[120] = 128;
	assign rom_real_data[121] = 99;
	assign rom_real_data[122] = 25;
	assign rom_real_data[123] = -60;
	assign rom_real_data[124] = -118;
	assign rom_real_data[125] = -122;
	assign rom_real_data[126] = -71;
	assign rom_real_data[127] = 13;
	assign rom_real_data[128] = 128;
	assign rom_real_data[129] = 128;
	assign rom_real_data[130] = 128;
	assign rom_real_data[131] = 128;
	assign rom_real_data[132] = 128;
	assign rom_real_data[133] = 128;
	assign rom_real_data[134] = 128;
	assign rom_real_data[135] = 128;
	assign rom_real_data[136] = 128;
	assign rom_real_data[137] = 118;
	assign rom_real_data[138] = 91;
	assign rom_real_data[139] = 49;
	assign rom_real_data[140] = 0;
	assign rom_real_data[141] = -49;
	assign rom_real_data[142] = -91;
	assign rom_real_data[143] = -118;
	assign rom_real_data[144] = 128;
	assign rom_real_data[145] = 126;
	assign rom_real_data[146] = 118;
	assign rom_real_data[147] = 106;
	assign rom_real_data[148] = 91;
	assign rom_real_data[149] = 71;
	assign rom_real_data[150] = 49;
	assign rom_real_data[151] = 25;
	assign rom_real_data[152] = 128;
	assign rom_real_data[153] = 106;
	assign rom_real_data[154] = 49;
	assign rom_real_data[155] = -25;
	assign rom_real_data[156] = -91;
	assign rom_real_data[157] = -126;
	assign rom_real_data[158] = -118;
	assign rom_real_data[159] = -71;
	assign rom_real_data[160] = 128;
	assign rom_real_data[161] = 127;
	assign rom_real_data[162] = 126;
	assign rom_real_data[163] = 122;
	assign rom_real_data[164] = 118;
	assign rom_real_data[165] = 113;
	assign rom_real_data[166] = 106;
	assign rom_real_data[167] = 99;
	assign rom_real_data[168] = 128;
	assign rom_real_data[169] = 113;
	assign rom_real_data[170] = 71;
	assign rom_real_data[171] = 13;
	assign rom_real_data[172] = -49;
	assign rom_real_data[173] = -99;
	assign rom_real_data[174] = -126;
	assign rom_real_data[175] = -122;
	assign rom_real_data[176] = 128;
	assign rom_real_data[177] = 122;
	assign rom_real_data[178] = 106;
	assign rom_real_data[179] = 81;
	assign rom_real_data[180] = 49;
	assign rom_real_data[181] = 13;
	assign rom_real_data[182] = -25;
	assign rom_real_data[183] = -60;
	assign rom_real_data[184] = 128;
	assign rom_real_data[185] = 99;
	assign rom_real_data[186] = 25;
	assign rom_real_data[187] = -60;
	assign rom_real_data[188] = -118;
	assign rom_real_data[189] = -122;
	assign rom_real_data[190] = -71;
	assign rom_real_data[191] = 13;
	assign rom_real_data[192] = 128;
	assign rom_real_data[193] = 128;
	assign rom_real_data[194] = 128;
	assign rom_real_data[195] = 128;
	assign rom_real_data[196] = 128;
	assign rom_real_data[197] = 128;
	assign rom_real_data[198] = 128;
	assign rom_real_data[199] = 128;
	assign rom_real_data[200] = 128;
	assign rom_real_data[201] = 118;
	assign rom_real_data[202] = 91;
	assign rom_real_data[203] = 49;
	assign rom_real_data[204] = 0;
	assign rom_real_data[205] = -49;
	assign rom_real_data[206] = -91;
	assign rom_real_data[207] = -118;
	assign rom_real_data[208] = 128;
	assign rom_real_data[209] = 126;
	assign rom_real_data[210] = 118;
	assign rom_real_data[211] = 106;
	assign rom_real_data[212] = 91;
	assign rom_real_data[213] = 71;
	assign rom_real_data[214] = 49;
	assign rom_real_data[215] = 25;
	assign rom_real_data[216] = 128;
	assign rom_real_data[217] = 106;
	assign rom_real_data[218] = 49;
	assign rom_real_data[219] = -25;
	assign rom_real_data[220] = -91;
	assign rom_real_data[221] = -126;
	assign rom_real_data[222] = -118;
	assign rom_real_data[223] = -71;
	assign rom_real_data[224] = 128;
	assign rom_real_data[225] = 127;
	assign rom_real_data[226] = 126;
	assign rom_real_data[227] = 122;
	assign rom_real_data[228] = 118;
	assign rom_real_data[229] = 113;
	assign rom_real_data[230] = 106;
	assign rom_real_data[231] = 99;
	assign rom_real_data[232] = 128;
	assign rom_real_data[233] = 113;
	assign rom_real_data[234] = 71;
	assign rom_real_data[235] = 13;
	assign rom_real_data[236] = -49;
	assign rom_real_data[237] = -99;
	assign rom_real_data[238] = -126;
	assign rom_real_data[239] = -122;
	assign rom_real_data[240] = 128;
	assign rom_real_data[241] = 122;
	assign rom_real_data[242] = 106;
	assign rom_real_data[243] = 81;
	assign rom_real_data[244] = 49;
	assign rom_real_data[245] = 13;
	assign rom_real_data[246] = -25;
	assign rom_real_data[247] = -60;
	assign rom_real_data[248] = 128;
	assign rom_real_data[249] = 99;
	assign rom_real_data[250] = 25;
	assign rom_real_data[251] = -60;
	assign rom_real_data[252] = -118;
	assign rom_real_data[253] = -122;
	assign rom_real_data[254] = -71;
	assign rom_real_data[255] = 13;
	assign rom_real_data[256] = 128;
	assign rom_real_data[257] = 128;
	assign rom_real_data[258] = 128;
	assign rom_real_data[259] = 128;
	assign rom_real_data[260] = 128;
	assign rom_real_data[261] = 128;
	assign rom_real_data[262] = 128;
	assign rom_real_data[263] = 128;
	assign rom_real_data[264] = 128;
	assign rom_real_data[265] = 118;
	assign rom_real_data[266] = 91;
	assign rom_real_data[267] = 49;
	assign rom_real_data[268] = 0;
	assign rom_real_data[269] = -49;
	assign rom_real_data[270] = -91;
	assign rom_real_data[271] = -118;
	assign rom_real_data[272] = 128;
	assign rom_real_data[273] = 126;
	assign rom_real_data[274] = 118;
	assign rom_real_data[275] = 106;
	assign rom_real_data[276] = 91;
	assign rom_real_data[277] = 71;
	assign rom_real_data[278] = 49;
	assign rom_real_data[279] = 25;
	assign rom_real_data[280] = 128;
	assign rom_real_data[281] = 106;
	assign rom_real_data[282] = 49;
	assign rom_real_data[283] = -25;
	assign rom_real_data[284] = -91;
	assign rom_real_data[285] = -126;
	assign rom_real_data[286] = -118;
	assign rom_real_data[287] = -71;
	assign rom_real_data[288] = 128;
	assign rom_real_data[289] = 127;
	assign rom_real_data[290] = 126;
	assign rom_real_data[291] = 122;
	assign rom_real_data[292] = 118;
	assign rom_real_data[293] = 113;
	assign rom_real_data[294] = 106;
	assign rom_real_data[295] = 99;
	assign rom_real_data[296] = 128;
	assign rom_real_data[297] = 113;
	assign rom_real_data[298] = 71;
	assign rom_real_data[299] = 13;
	assign rom_real_data[300] = -49;
	assign rom_real_data[301] = -99;
	assign rom_real_data[302] = -126;
	assign rom_real_data[303] = -122;
	assign rom_real_data[304] = 128;
	assign rom_real_data[305] = 122;
	assign rom_real_data[306] = 106;
	assign rom_real_data[307] = 81;
	assign rom_real_data[308] = 49;
	assign rom_real_data[309] = 13;
	assign rom_real_data[310] = -25;
	assign rom_real_data[311] = -60;
	assign rom_real_data[312] = 128;
	assign rom_real_data[313] = 99;
	assign rom_real_data[314] = 25;
	assign rom_real_data[315] = -60;
	assign rom_real_data[316] = -118;
	assign rom_real_data[317] = -122;
	assign rom_real_data[318] = -71;
	assign rom_real_data[319] = 13;
	assign rom_real_data[320] = 128;
	assign rom_real_data[321] = 128;
	assign rom_real_data[322] = 128;
	assign rom_real_data[323] = 128;
	assign rom_real_data[324] = 128;
	assign rom_real_data[325] = 128;
	assign rom_real_data[326] = 128;
	assign rom_real_data[327] = 128;
	assign rom_real_data[328] = 128;
	assign rom_real_data[329] = 118;
	assign rom_real_data[330] = 91;
	assign rom_real_data[331] = 49;
	assign rom_real_data[332] = 0;
	assign rom_real_data[333] = -49;
	assign rom_real_data[334] = -91;
	assign rom_real_data[335] = -118;
	assign rom_real_data[336] = 128;
	assign rom_real_data[337] = 126;
	assign rom_real_data[338] = 118;
	assign rom_real_data[339] = 106;
	assign rom_real_data[340] = 91;
	assign rom_real_data[341] = 71;
	assign rom_real_data[342] = 49;
	assign rom_real_data[343] = 25;
	assign rom_real_data[344] = 128;
	assign rom_real_data[345] = 106;
	assign rom_real_data[346] = 49;
	assign rom_real_data[347] = -25;
	assign rom_real_data[348] = -91;
	assign rom_real_data[349] = -126;
	assign rom_real_data[350] = -118;
	assign rom_real_data[351] = -71;
	assign rom_real_data[352] = 128;
	assign rom_real_data[353] = 127;
	assign rom_real_data[354] = 126;
	assign rom_real_data[355] = 122;
	assign rom_real_data[356] = 118;
	assign rom_real_data[357] = 113;
	assign rom_real_data[358] = 106;
	assign rom_real_data[359] = 99;
	assign rom_real_data[360] = 128;
	assign rom_real_data[361] = 113;
	assign rom_real_data[362] = 71;
	assign rom_real_data[363] = 13;
	assign rom_real_data[364] = -49;
	assign rom_real_data[365] = -99;
	assign rom_real_data[366] = -126;
	assign rom_real_data[367] = -122;
	assign rom_real_data[368] = 128;
	assign rom_real_data[369] = 122;
	assign rom_real_data[370] = 106;
	assign rom_real_data[371] = 81;
	assign rom_real_data[372] = 49;
	assign rom_real_data[373] = 13;
	assign rom_real_data[374] = -25;
	assign rom_real_data[375] = -60;
	assign rom_real_data[376] = 128;
	assign rom_real_data[377] = 99;
	assign rom_real_data[378] = 25;
	assign rom_real_data[379] = -60;
	assign rom_real_data[380] = -118;
	assign rom_real_data[381] = -122;
	assign rom_real_data[382] = -71;
	assign rom_real_data[383] = 13;
	assign rom_real_data[384] = 128;
	assign rom_real_data[385] = 128;
	assign rom_real_data[386] = 128;
	assign rom_real_data[387] = 128;
	assign rom_real_data[388] = 128;
	assign rom_real_data[389] = 128;
	assign rom_real_data[390] = 128;
	assign rom_real_data[391] = 128;
	assign rom_real_data[392] = 128;
	assign rom_real_data[393] = 118;
	assign rom_real_data[394] = 91;
	assign rom_real_data[395] = 49;
	assign rom_real_data[396] = 0;
	assign rom_real_data[397] = -49;
	assign rom_real_data[398] = -91;
	assign rom_real_data[399] = -118;
	assign rom_real_data[400] = 128;
	assign rom_real_data[401] = 126;
	assign rom_real_data[402] = 118;
	assign rom_real_data[403] = 106;
	assign rom_real_data[404] = 91;
	assign rom_real_data[405] = 71;
	assign rom_real_data[406] = 49;
	assign rom_real_data[407] = 25;
	assign rom_real_data[408] = 128;
	assign rom_real_data[409] = 106;
	assign rom_real_data[410] = 49;
	assign rom_real_data[411] = -25;
	assign rom_real_data[412] = -91;
	assign rom_real_data[413] = -126;
	assign rom_real_data[414] = -118;
	assign rom_real_data[415] = -71;
	assign rom_real_data[416] = 128;
	assign rom_real_data[417] = 127;
	assign rom_real_data[418] = 126;
	assign rom_real_data[419] = 122;
	assign rom_real_data[420] = 118;
	assign rom_real_data[421] = 113;
	assign rom_real_data[422] = 106;
	assign rom_real_data[423] = 99;
	assign rom_real_data[424] = 128;
	assign rom_real_data[425] = 113;
	assign rom_real_data[426] = 71;
	assign rom_real_data[427] = 13;
	assign rom_real_data[428] = -49;
	assign rom_real_data[429] = -99;
	assign rom_real_data[430] = -126;
	assign rom_real_data[431] = -122;
	assign rom_real_data[432] = 128;
	assign rom_real_data[433] = 122;
	assign rom_real_data[434] = 106;
	assign rom_real_data[435] = 81;
	assign rom_real_data[436] = 49;
	assign rom_real_data[437] = 13;
	assign rom_real_data[438] = -25;
	assign rom_real_data[439] = -60;
	assign rom_real_data[440] = 128;
	assign rom_real_data[441] = 99;
	assign rom_real_data[442] = 25;
	assign rom_real_data[443] = -60;
	assign rom_real_data[444] = -118;
	assign rom_real_data[445] = -122;
	assign rom_real_data[446] = -71;
	assign rom_real_data[447] = 13;
	assign rom_real_data[448] = 128;
	assign rom_real_data[449] = 128;
	assign rom_real_data[450] = 128;
	assign rom_real_data[451] = 128;
	assign rom_real_data[452] = 128;
	assign rom_real_data[453] = 128;
	assign rom_real_data[454] = 128;
	assign rom_real_data[455] = 128;
	assign rom_real_data[456] = 128;
	assign rom_real_data[457] = 118;
	assign rom_real_data[458] = 91;
	assign rom_real_data[459] = 49;
	assign rom_real_data[460] = 0;
	assign rom_real_data[461] = -49;
	assign rom_real_data[462] = -91;
	assign rom_real_data[463] = -118;
	assign rom_real_data[464] = 128;
	assign rom_real_data[465] = 126;
	assign rom_real_data[466] = 118;
	assign rom_real_data[467] = 106;
	assign rom_real_data[468] = 91;
	assign rom_real_data[469] = 71;
	assign rom_real_data[470] = 49;
	assign rom_real_data[471] = 25;
	assign rom_real_data[472] = 128;
	assign rom_real_data[473] = 106;
	assign rom_real_data[474] = 49;
	assign rom_real_data[475] = -25;
	assign rom_real_data[476] = -91;
	assign rom_real_data[477] = -126;
	assign rom_real_data[478] = -118;
	assign rom_real_data[479] = -71;
	assign rom_real_data[480] = 128;
	assign rom_real_data[481] = 127;
	assign rom_real_data[482] = 126;
	assign rom_real_data[483] = 122;
	assign rom_real_data[484] = 118;
	assign rom_real_data[485] = 113;
	assign rom_real_data[486] = 106;
	assign rom_real_data[487] = 99;
	assign rom_real_data[488] = 128;
	assign rom_real_data[489] = 113;
	assign rom_real_data[490] = 71;
	assign rom_real_data[491] = 13;
	assign rom_real_data[492] = -49;
	assign rom_real_data[493] = -99;
	assign rom_real_data[494] = -126;
	assign rom_real_data[495] = -122;
	assign rom_real_data[496] = 128;
	assign rom_real_data[497] = 122;
	assign rom_real_data[498] = 106;
	assign rom_real_data[499] = 81;
	assign rom_real_data[500] = 49;
	assign rom_real_data[501] = 13;
	assign rom_real_data[502] = -25;
	assign rom_real_data[503] = -60;
	assign rom_real_data[504] = 128;
	assign rom_real_data[505] = 99;
	assign rom_real_data[506] = 25;
	assign rom_real_data[507] = -60;
	assign rom_real_data[508] = -118;
	assign rom_real_data[509] = -122;
	assign rom_real_data[510] = -71;
	assign rom_real_data[511] = 13;


	assign rom_imag_data[0]   = 0;
	assign rom_imag_data[1]   = 0;
	assign rom_imag_data[2]   = 0;
	assign rom_imag_data[3]   = 0;
	assign rom_imag_data[4]   = 0;
	assign rom_imag_data[5]   = 0;
	assign rom_imag_data[6]   = 0;
	assign rom_imag_data[7]   = 0;
	assign rom_imag_data[8]   = 0;
	assign rom_imag_data[9]   = -49;
	assign rom_imag_data[10]  = -91;
	assign rom_imag_data[11]  = -118;
	assign rom_imag_data[12]  = -128;
	assign rom_imag_data[13]  = -118;
	assign rom_imag_data[14]  = -91;
	assign rom_imag_data[15]  = -49;
	assign rom_imag_data[16]  = 0;
	assign rom_imag_data[17]  = -25;
	assign rom_imag_data[18]  = -49;
	assign rom_imag_data[19]  = -71;
	assign rom_imag_data[20]  = -91;
	assign rom_imag_data[21]  = -106;
	assign rom_imag_data[22]  = -118;
	assign rom_imag_data[23]  = -126;
	assign rom_imag_data[24]  = 0;
	assign rom_imag_data[25]  = -71;
	assign rom_imag_data[26]  = -118;
	assign rom_imag_data[27]  = -126;
	assign rom_imag_data[28]  = -91;
	assign rom_imag_data[29]  = -25;
	assign rom_imag_data[30]  = 49;
	assign rom_imag_data[31]  = 106;
	assign rom_imag_data[32]  = 0;
	assign rom_imag_data[33]  = -13;
	assign rom_imag_data[34]  = -25;
	assign rom_imag_data[35]  = -37;
	assign rom_imag_data[36]  = -49;
	assign rom_imag_data[37]  = -60;
	assign rom_imag_data[38]  = -71;
	assign rom_imag_data[39]  = -81;
	assign rom_imag_data[40]  = 0;
	assign rom_imag_data[41]  = -60;
	assign rom_imag_data[42]  = -106;
	assign rom_imag_data[43]  = -127;
	assign rom_imag_data[44]  = -118;
	assign rom_imag_data[45]  = -81;
	assign rom_imag_data[46]  = -25;
	assign rom_imag_data[47]  = 37;
	assign rom_imag_data[48]  = 0;
	assign rom_imag_data[49]  = -37;
	assign rom_imag_data[50]  = -71;
	assign rom_imag_data[51]  = -99;
	assign rom_imag_data[52]  = -118;
	assign rom_imag_data[53]  = -127;
	assign rom_imag_data[54]  = -126;
	assign rom_imag_data[55]  = -113;
	assign rom_imag_data[56]  = 0;
	assign rom_imag_data[57]  = -81;
	assign rom_imag_data[58]  = -126;
	assign rom_imag_data[59]  = -113;
	assign rom_imag_data[60]  = -49;
	assign rom_imag_data[61]  = 37;
	assign rom_imag_data[62]  = 106;
	assign rom_imag_data[63]  = 127;
	assign rom_imag_data[64]  = 0;
	assign rom_imag_data[65]  = 0;
	assign rom_imag_data[66]  = 0;
	assign rom_imag_data[67]  = 0;
	assign rom_imag_data[68]  = 0;
	assign rom_imag_data[69]  = 0;
	assign rom_imag_data[70]  = 0;
	assign rom_imag_data[71]  = 0;
	assign rom_imag_data[72]  = 0;
	assign rom_imag_data[73]  = -49;
	assign rom_imag_data[74]  = -91;
	assign rom_imag_data[75]  = -118;
	assign rom_imag_data[76]  = -128;
	assign rom_imag_data[77]  = -118;
	assign rom_imag_data[78]  = -91;
	assign rom_imag_data[79]  = -49;
	assign rom_imag_data[80]  = 0;
	assign rom_imag_data[81]  = -25;
	assign rom_imag_data[82]  = -49;
	assign rom_imag_data[83]  = -71;
	assign rom_imag_data[84]  = -91;
	assign rom_imag_data[85]  = -106;
	assign rom_imag_data[86]  = -118;
	assign rom_imag_data[87]  = -126;
	assign rom_imag_data[88]  = 0;
	assign rom_imag_data[89]  = -71;
	assign rom_imag_data[90]  = -118;
	assign rom_imag_data[91]  = -126;
	assign rom_imag_data[92]  = -91;
	assign rom_imag_data[93]  = -25;
	assign rom_imag_data[94]  = 49;
	assign rom_imag_data[95]  = 106;
	assign rom_imag_data[96]  = 0;
	assign rom_imag_data[97]  = -13;
	assign rom_imag_data[98]  = -25;
	assign rom_imag_data[99]  = -37;
	assign rom_imag_data[100] = -49;
	assign rom_imag_data[101] = -60;
	assign rom_imag_data[102] = -71;
	assign rom_imag_data[103] = -81;
	assign rom_imag_data[104] = 0;
	assign rom_imag_data[105] = -60;
	assign rom_imag_data[106] = -106;
	assign rom_imag_data[107] = -127;
	assign rom_imag_data[108] = -118;
	assign rom_imag_data[109] = -81;
	assign rom_imag_data[110] = -25;
	assign rom_imag_data[111] = 37;
	assign rom_imag_data[112] = 0;
	assign rom_imag_data[113] = -37;
	assign rom_imag_data[114] = -71;
	assign rom_imag_data[115] = -99;
	assign rom_imag_data[116] = -118;
	assign rom_imag_data[117] = -127;
	assign rom_imag_data[118] = -126;
	assign rom_imag_data[119] = -113;
	assign rom_imag_data[120] = 0;
	assign rom_imag_data[121] = -81;
	assign rom_imag_data[122] = -126;
	assign rom_imag_data[123] = -113;
	assign rom_imag_data[124] = -49;
	assign rom_imag_data[125] = 37;
	assign rom_imag_data[126] = 106;
	assign rom_imag_data[127] = 127;
	assign rom_imag_data[128] = 0;
	assign rom_imag_data[129] = 0;
	assign rom_imag_data[130] = 0;
	assign rom_imag_data[131] = 0;
	assign rom_imag_data[132] = 0;
	assign rom_imag_data[133] = 0;
	assign rom_imag_data[134] = 0;
	assign rom_imag_data[135] = 0;
	assign rom_imag_data[136] = 0;
	assign rom_imag_data[137] = -49;
	assign rom_imag_data[138] = -91;
	assign rom_imag_data[139] = -118;
	assign rom_imag_data[140] = -128;
	assign rom_imag_data[141] = -118;
	assign rom_imag_data[142] = -91;
	assign rom_imag_data[143] = -49;
	assign rom_imag_data[144] = 0;
	assign rom_imag_data[145] = -25;
	assign rom_imag_data[146] = -49;
	assign rom_imag_data[147] = -71;
	assign rom_imag_data[148] = -91;
	assign rom_imag_data[149] = -106;
	assign rom_imag_data[150] = -118;
	assign rom_imag_data[151] = -126;
	assign rom_imag_data[152] = 0;
	assign rom_imag_data[153] = -71;
	assign rom_imag_data[154] = -118;
	assign rom_imag_data[155] = -126;
	assign rom_imag_data[156] = -91;
	assign rom_imag_data[157] = -25;
	assign rom_imag_data[158] = 49;
	assign rom_imag_data[159] = 106;
	assign rom_imag_data[160] = 0;
	assign rom_imag_data[161] = -13;
	assign rom_imag_data[162] = -25;
	assign rom_imag_data[163] = -37;
	assign rom_imag_data[164] = -49;
	assign rom_imag_data[165] = -60;
	assign rom_imag_data[166] = -71;
	assign rom_imag_data[167] = -81;
	assign rom_imag_data[168] = 0;
	assign rom_imag_data[169] = -60;
	assign rom_imag_data[170] = -106;
	assign rom_imag_data[171] = -127;
	assign rom_imag_data[172] = -118;
	assign rom_imag_data[173] = -81;
	assign rom_imag_data[174] = -25;
	assign rom_imag_data[175] = 37;
	assign rom_imag_data[176] = 0;
	assign rom_imag_data[177] = -37;
	assign rom_imag_data[178] = -71;
	assign rom_imag_data[179] = -99;
	assign rom_imag_data[180] = -118;
	assign rom_imag_data[181] = -127;
	assign rom_imag_data[182] = -126;
	assign rom_imag_data[183] = -113;
	assign rom_imag_data[184] = 0;
	assign rom_imag_data[185] = -81;
	assign rom_imag_data[186] = -126;
	assign rom_imag_data[187] = -113;
	assign rom_imag_data[188] = -49;
	assign rom_imag_data[189] = 37;
	assign rom_imag_data[190] = 106;
	assign rom_imag_data[191] = 127;
	assign rom_imag_data[192] = 0;
	assign rom_imag_data[193] = 0;
	assign rom_imag_data[194] = 0;
	assign rom_imag_data[195] = 0;
	assign rom_imag_data[196] = 0;
	assign rom_imag_data[197] = 0;
	assign rom_imag_data[198] = 0;
	assign rom_imag_data[199] = 0;
	assign rom_imag_data[200] = 0;
	assign rom_imag_data[201] = -49;
	assign rom_imag_data[202] = -91;
	assign rom_imag_data[203] = -118;
	assign rom_imag_data[204] = -128;
	assign rom_imag_data[205] = -118;
	assign rom_imag_data[206] = -91;
	assign rom_imag_data[207] = -49;
	assign rom_imag_data[208] = 0;
	assign rom_imag_data[209] = -25;
	assign rom_imag_data[210] = -49;
	assign rom_imag_data[211] = -71;
	assign rom_imag_data[212] = -91;
	assign rom_imag_data[213] = -106;
	assign rom_imag_data[214] = -118;
	assign rom_imag_data[215] = -126;
	assign rom_imag_data[216] = 0;
	assign rom_imag_data[217] = -71;
	assign rom_imag_data[218] = -118;
	assign rom_imag_data[219] = -126;
	assign rom_imag_data[220] = -91;
	assign rom_imag_data[221] = -25;
	assign rom_imag_data[222] = 49;
	assign rom_imag_data[223] = 106;
	assign rom_imag_data[224] = 0;
	assign rom_imag_data[225] = -13;
	assign rom_imag_data[226] = -25;
	assign rom_imag_data[227] = -37;
	assign rom_imag_data[228] = -49;
	assign rom_imag_data[229] = -60;
	assign rom_imag_data[230] = -71;
	assign rom_imag_data[231] = -81;
	assign rom_imag_data[232] = 0;
	assign rom_imag_data[233] = -60;
	assign rom_imag_data[234] = -106;
	assign rom_imag_data[235] = -127;
	assign rom_imag_data[236] = -118;
	assign rom_imag_data[237] = -81;
	assign rom_imag_data[238] = -25;
	assign rom_imag_data[239] = 37;
	assign rom_imag_data[240] = 0;
	assign rom_imag_data[241] = -37;
	assign rom_imag_data[242] = -71;
	assign rom_imag_data[243] = -99;
	assign rom_imag_data[244] = -118;
	assign rom_imag_data[245] = -127;
	assign rom_imag_data[246] = -126;
	assign rom_imag_data[247] = -113;
	assign rom_imag_data[248] = 0;
	assign rom_imag_data[249] = -81;
	assign rom_imag_data[250] = -126;
	assign rom_imag_data[251] = -113;
	assign rom_imag_data[252] = -49;
	assign rom_imag_data[253] = 37;
	assign rom_imag_data[254] = 106;
	assign rom_imag_data[255] = 127;
	assign rom_imag_data[256] = 0;
	assign rom_imag_data[257] = 0;
	assign rom_imag_data[258] = 0;
	assign rom_imag_data[259] = 0;
	assign rom_imag_data[260] = 0;
	assign rom_imag_data[261] = 0;
	assign rom_imag_data[262] = 0;
	assign rom_imag_data[263] = 0;
	assign rom_imag_data[264] = 0;
	assign rom_imag_data[265] = -49;
	assign rom_imag_data[266] = -91;
	assign rom_imag_data[267] = -118;
	assign rom_imag_data[268] = -128;
	assign rom_imag_data[269] = -118;
	assign rom_imag_data[270] = -91;
	assign rom_imag_data[271] = -49;
	assign rom_imag_data[272] = 0;
	assign rom_imag_data[273] = -25;
	assign rom_imag_data[274] = -49;
	assign rom_imag_data[275] = -71;
	assign rom_imag_data[276] = -91;
	assign rom_imag_data[277] = -106;
	assign rom_imag_data[278] = -118;
	assign rom_imag_data[279] = -126;
	assign rom_imag_data[280] = 0;
	assign rom_imag_data[281] = -71;
	assign rom_imag_data[282] = -118;
	assign rom_imag_data[283] = -126;
	assign rom_imag_data[284] = -91;
	assign rom_imag_data[285] = -25;
	assign rom_imag_data[286] = 49;
	assign rom_imag_data[287] = 106;
	assign rom_imag_data[288] = 0;
	assign rom_imag_data[289] = -13;
	assign rom_imag_data[290] = -25;
	assign rom_imag_data[291] = -37;
	assign rom_imag_data[292] = -49;
	assign rom_imag_data[293] = -60;
	assign rom_imag_data[294] = -71;
	assign rom_imag_data[295] = -81;
	assign rom_imag_data[296] = 0;
	assign rom_imag_data[297] = -60;
	assign rom_imag_data[298] = -106;
	assign rom_imag_data[299] = -127;
	assign rom_imag_data[300] = -118;
	assign rom_imag_data[301] = -81;
	assign rom_imag_data[302] = -25;
	assign rom_imag_data[303] = 37;
	assign rom_imag_data[304] = 0;
	assign rom_imag_data[305] = -37;
	assign rom_imag_data[306] = -71;
	assign rom_imag_data[307] = -99;
	assign rom_imag_data[308] = -118;
	assign rom_imag_data[309] = -127;
	assign rom_imag_data[310] = -126;
	assign rom_imag_data[311] = -113;
	assign rom_imag_data[312] = 0;
	assign rom_imag_data[313] = -81;
	assign rom_imag_data[314] = -126;
	assign rom_imag_data[315] = -113;
	assign rom_imag_data[316] = -49;
	assign rom_imag_data[317] = 37;
	assign rom_imag_data[318] = 106;
	assign rom_imag_data[319] = 127;
	assign rom_imag_data[320] = 0;
	assign rom_imag_data[321] = 0;
	assign rom_imag_data[322] = 0;
	assign rom_imag_data[323] = 0;
	assign rom_imag_data[324] = 0;
	assign rom_imag_data[325] = 0;
	assign rom_imag_data[326] = 0;
	assign rom_imag_data[327] = 0;
	assign rom_imag_data[328] = 0;
	assign rom_imag_data[329] = -49;
	assign rom_imag_data[330] = -91;
	assign rom_imag_data[331] = -118;
	assign rom_imag_data[332] = -128;
	assign rom_imag_data[333] = -118;
	assign rom_imag_data[334] = -91;
	assign rom_imag_data[335] = -49;
	assign rom_imag_data[336] = 0;
	assign rom_imag_data[337] = -25;
	assign rom_imag_data[338] = -49;
	assign rom_imag_data[339] = -71;
	assign rom_imag_data[340] = -91;
	assign rom_imag_data[341] = -106;
	assign rom_imag_data[342] = -118;
	assign rom_imag_data[343] = -126;
	assign rom_imag_data[344] = 0;
	assign rom_imag_data[345] = -71;
	assign rom_imag_data[346] = -118;
	assign rom_imag_data[347] = -126;
	assign rom_imag_data[348] = -91;
	assign rom_imag_data[349] = -25;
	assign rom_imag_data[350] = 49;
	assign rom_imag_data[351] = 106;
	assign rom_imag_data[352] = 0;
	assign rom_imag_data[353] = -13;
	assign rom_imag_data[354] = -25;
	assign rom_imag_data[355] = -37;
	assign rom_imag_data[356] = -49;
	assign rom_imag_data[357] = -60;
	assign rom_imag_data[358] = -71;
	assign rom_imag_data[359] = -81;
	assign rom_imag_data[360] = 0;
	assign rom_imag_data[361] = -60;
	assign rom_imag_data[362] = -106;
	assign rom_imag_data[363] = -127;
	assign rom_imag_data[364] = -118;
	assign rom_imag_data[365] = -81;
	assign rom_imag_data[366] = -25;
	assign rom_imag_data[367] = 37;
	assign rom_imag_data[368] = 0;
	assign rom_imag_data[369] = -37;
	assign rom_imag_data[370] = -71;
	assign rom_imag_data[371] = -99;
	assign rom_imag_data[372] = -118;
	assign rom_imag_data[373] = -127;
	assign rom_imag_data[374] = -126;
	assign rom_imag_data[375] = -113;
	assign rom_imag_data[376] = 0;
	assign rom_imag_data[377] = -81;
	assign rom_imag_data[378] = -126;
	assign rom_imag_data[379] = -113;
	assign rom_imag_data[380] = -49;
	assign rom_imag_data[381] = 37;
	assign rom_imag_data[382] = 106;
	assign rom_imag_data[383] = 127;
	assign rom_imag_data[384] = 0;
	assign rom_imag_data[385] = 0;
	assign rom_imag_data[386] = 0;
	assign rom_imag_data[387] = 0;
	assign rom_imag_data[388] = 0;
	assign rom_imag_data[389] = 0;
	assign rom_imag_data[390] = 0;
	assign rom_imag_data[391] = 0;
	assign rom_imag_data[392] = 0;
	assign rom_imag_data[393] = -49;
	assign rom_imag_data[394] = -91;
	assign rom_imag_data[395] = -118;
	assign rom_imag_data[396] = -128;
	assign rom_imag_data[397] = -118;
	assign rom_imag_data[398] = -91;
	assign rom_imag_data[399] = -49;
	assign rom_imag_data[400] = 0;
	assign rom_imag_data[401] = -25;
	assign rom_imag_data[402] = -49;
	assign rom_imag_data[403] = -71;
	assign rom_imag_data[404] = -91;
	assign rom_imag_data[405] = -106;
	assign rom_imag_data[406] = -118;
	assign rom_imag_data[407] = -126;
	assign rom_imag_data[408] = 0;
	assign rom_imag_data[409] = -71;
	assign rom_imag_data[410] = -118;
	assign rom_imag_data[411] = -126;
	assign rom_imag_data[412] = -91;
	assign rom_imag_data[413] = -25;
	assign rom_imag_data[414] = 49;
	assign rom_imag_data[415] = 106;
	assign rom_imag_data[416] = 0;
	assign rom_imag_data[417] = -13;
	assign rom_imag_data[418] = -25;
	assign rom_imag_data[419] = -37;
	assign rom_imag_data[420] = -49;
	assign rom_imag_data[421] = -60;
	assign rom_imag_data[422] = -71;
	assign rom_imag_data[423] = -81;
	assign rom_imag_data[424] = 0;
	assign rom_imag_data[425] = -60;
	assign rom_imag_data[426] = -106;
	assign rom_imag_data[427] = -127;
	assign rom_imag_data[428] = -118;
	assign rom_imag_data[429] = -81;
	assign rom_imag_data[430] = -25;
	assign rom_imag_data[431] = 37;
	assign rom_imag_data[432] = 0;
	assign rom_imag_data[433] = -37;
	assign rom_imag_data[434] = -71;
	assign rom_imag_data[435] = -99;
	assign rom_imag_data[436] = -118;
	assign rom_imag_data[437] = -127;
	assign rom_imag_data[438] = -126;
	assign rom_imag_data[439] = -113;
	assign rom_imag_data[440] = 0;
	assign rom_imag_data[441] = -81;
	assign rom_imag_data[442] = -126;
	assign rom_imag_data[443] = -113;
	assign rom_imag_data[444] = -49;
	assign rom_imag_data[445] = 37;
	assign rom_imag_data[446] = 106;
	assign rom_imag_data[447] = 127;
	assign rom_imag_data[448] = 0;
	assign rom_imag_data[449] = 0;
	assign rom_imag_data[450] = 0;
	assign rom_imag_data[451] = 0;
	assign rom_imag_data[452] = 0;
	assign rom_imag_data[453] = 0;
	assign rom_imag_data[454] = 0;
	assign rom_imag_data[455] = 0;
	assign rom_imag_data[456] = 0;
	assign rom_imag_data[457] = -49;
	assign rom_imag_data[458] = -91;
	assign rom_imag_data[459] = -118;
	assign rom_imag_data[460] = -128;
	assign rom_imag_data[461] = -118;
	assign rom_imag_data[462] = -91;
	assign rom_imag_data[463] = -49;
	assign rom_imag_data[464] = 0;
	assign rom_imag_data[465] = -25;
	assign rom_imag_data[466] = -49;
	assign rom_imag_data[467] = -71;
	assign rom_imag_data[468] = -91;
	assign rom_imag_data[469] = -106;
	assign rom_imag_data[470] = -118;
	assign rom_imag_data[471] = -126;
	assign rom_imag_data[472] = 0;
	assign rom_imag_data[473] = -71;
	assign rom_imag_data[474] = -118;
	assign rom_imag_data[475] = -126;
	assign rom_imag_data[476] = -91;
	assign rom_imag_data[477] = -25;
	assign rom_imag_data[478] = 49;
	assign rom_imag_data[479] = 106;
	assign rom_imag_data[480] = 0;
	assign rom_imag_data[481] = -13;
	assign rom_imag_data[482] = -25;
	assign rom_imag_data[483] = -37;
	assign rom_imag_data[484] = -49;
	assign rom_imag_data[485] = -60;
	assign rom_imag_data[486] = -71;
	assign rom_imag_data[487] = -81;
	assign rom_imag_data[488] = 0;
	assign rom_imag_data[489] = -60;
	assign rom_imag_data[490] = -106;
	assign rom_imag_data[491] = -127;
	assign rom_imag_data[492] = -118;
	assign rom_imag_data[493] = -81;
	assign rom_imag_data[494] = -25;
	assign rom_imag_data[495] = 37;
	assign rom_imag_data[496] = 0;
	assign rom_imag_data[497] = -37;
	assign rom_imag_data[498] = -71;
	assign rom_imag_data[499] = -99;
	assign rom_imag_data[500] = -118;
	assign rom_imag_data[501] = -127;
	assign rom_imag_data[502] = -126;
	assign rom_imag_data[503] = -113;
	assign rom_imag_data[504] = 0;
	assign rom_imag_data[505] = -81;
	assign rom_imag_data[506] = -126;
	assign rom_imag_data[507] = -113;
	assign rom_imag_data[508] = -49;
	assign rom_imag_data[509] = 37;
	assign rom_imag_data[510] = 106;
	assign rom_imag_data[511] = 127;

    
endmodule
